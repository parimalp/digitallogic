`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Module Name: xup_or3
//////////////////////////////////////////////////////////////////////////////////
module xup_or3 #(parameter DELAY = 3)(
    input wire a,
    input wire b,
    input wire c,
    output wire y
    );
    
    or #DELAY (y,a,b,c);
    
endmodule
