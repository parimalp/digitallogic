`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Module Name: xup_and3
//////////////////////////////////////////////////////////////////////////////////
module xup_and3 #(parameter DELAY=3)(
    input wire a,
    input wire b,
    input wire c,
    output wire y
    );
    
    and #DELAY (y,a,b,c);
    
endmodule
