`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Module Name: xup_or2
//////////////////////////////////////////////////////////////////////////////////
module xup_or2 #(parameter DELAY = 3)(
    input wire a,
    input wire b,
    output wire y
    );
    
    or #DELAY (y,a,b);
    
endmodule
